`include "defines.sv" 
module rom(
    input InstAddrBus pc_i,

    output InstBus    inst
);
always_comb begin
    unique case (pc_i)
        8'd0    : inst <= 32'b000000000000_00000_000_0000_0010011;
        8'd1    : inst <= 32'b000000001111_00001_000_00001_0010011;
        8'd2    : inst <= 32'b000000001111_00001_000_00010_0010011;
        8'd3    : inst <= 32'b0000000_00010_00001_000_00001_0110011;
        8'd4    : inst <= 32'b0000000_00010_00001_000_00001_0110011;
        8'd5    : inst <= 32'b0000000_00010_00001_000_00001_0110011;
        8'd6    : inst <= 32'b0000000_00010_00001_000_00001_0110011;
        8'd7    : inst <= 32'b0000000_00010_00001_000_00001_0110011;
        default : inst <= 32'b000000000000_00000_000_0000_0010011;
    endcase
end
endmodule
