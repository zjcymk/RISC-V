package pkg;
    typedef struct  {
    logic clk;
    logic rst_n;
} sys_t;
endpackage